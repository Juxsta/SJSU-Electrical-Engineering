module Majority_Circuit(
    input A,
    input B,
    input C,
    input D,
    output M,
    output U,
    output T
);
    assign  M = 

endmodule